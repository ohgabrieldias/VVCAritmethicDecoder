module add_4(
    input wire [7:0] in,
    output wire [7:0] out
);
    assign out = in + 4;
endmodule