module right_shift_5(
    input wire [8:0] in,
    output wire [8:0] out
);
    assign out = in >> 5;
endmodule
